`timescale 1ns/1ps

// src/pcpi_sha.v
// Simple PCPI coprocessor implementing Sigma0(rs1) = ROTR(rs1,2) ^ ROTR(rs1,13) ^ ROTR(rs1,22).
// Matches the standard picorv32 pcpi interface: (pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2) -> (pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready)

module pcpi_sha (
    input  wire        pcpi_valid,
    input  wire [31:0] pcpi_insn,
    input  wire [31:0] pcpi_rs1,
    input  wire [31:0] pcpi_rs2,

    output reg         pcpi_wr,
    output reg [31:0]  pcpi_rd,
    output reg         pcpi_wait,
    output reg         pcpi_ready
);

    // instruction fields
    wire [6:0] opcode = pcpi_insn[6:0];
    wire [2:0] funct3 = pcpi_insn[14:12];

    localparam [6:0] OPC_CUSTOM0 = 7'b0001011; // CUSTOM_0 opcode

    function [31:0] rotr;
        input [31:0] x;
        input integer n;
        begin
            rotr = (x >> n) | (x << (32-n));
        end
    endfunction

    always @(*) begin
        pcpi_wr    = 1'b0;
        pcpi_rd    = 32'b0;
        pcpi_wait  = 1'b0;
        pcpi_ready = 1'b0;

        if (pcpi_valid) begin
            if ((opcode == OPC_CUSTOM0) && (funct3 == 3'b000)) begin
                pcpi_rd    = rotr(pcpi_rs1, 2) ^ rotr(pcpi_rs1, 13) ^ rotr(pcpi_rs1, 22);
                pcpi_wr    = 1'b1;
                pcpi_ready = 1'b1; // combinational ready
            end
        end
    end

endmodule
